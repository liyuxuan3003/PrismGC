module clk_200k( );



endmodule
