module clk1000HZ( );



endmodule
