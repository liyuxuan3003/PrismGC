`protect begin_protected
`protect version = 1
`protect encrypt_agent = "Anlogic"
`protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-002"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`protect key_block
QNadfMIDUn13TN6mqrK6CCwIDXvgNdUlFCpNp7x26cAfj6mPtUYrzsdyDlswD7Y4
bdUW2jxJK6XTpG4hSw42qwuWFZnMhVhFvqHFFmQDHAk1oKIDUHSzmliyDc05OLyu
7ofz78RnaasBna0CYAYlNd0cguqIB0zgkRbCfCFwCLc=
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`protect key_block
eAevTaLd62PHmOCX2kwDIs8Bs2Y1MkOFDf/0g0THDqhtvoi8s0cHqS+x4q04zsye
AdWvGVkk90OIi/glYGsyJMKrkzdeJJ6gXeOjqJGebHunE4Vixm4fZW7NLwfZfew3
Q4jEL95iTtVTOsWNYxFoJVm07Z/UEEy5mdxY+QnVRXJdSnwdsENJyXThSgAmL2PI
6uZ/YoJGi8ZRgtU6mrBhaCYtLyP8GmwRcxuGx/Qpy3z7rHh8fGgwmSfaVNtLSNvE
Z7yTwKKpwY3/OrUL6z8z/IXiyIqr3HaPZSN9Kz/0rvIme9wiijrCmeTNwzsWatSU
U+qO0TCo+FqWMfILKFR/Ag==
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`protect key_block
nRvoGpO5t+qt3hsG5A82aBgwgS3x9ZqDCgr3vQ0uIaaaDg/yTSIgfvEcaqVm9bMS
OiZ0kUcvQi29w7viwag2EoXbE58aZ5JDRm4L8nPCY0pfP9dphCnpmQMuXpp+EYRa
W6uiXnudrHcYgwIcX9aIs9Kc+bRQORksJutI0JTJxJM=
`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`protect key_block
d1tEbXyaZ5Fyn/5h2d57ySDaYPGFaY3i6j8qeL4gNIGVMUj0AgvPeekdiEiRZWKv
hqadidae/aEWMN3yRm7T1M7QWO7dUtNawXNmCp6gVdBKZwpT8oMhuJspvraz+aTE
VBMjrZVdgD+khbI5PURdQckQ6Bcf100Vs7tvvOPFxzYDOr47k+SRllpxj5lXo2jo
T9kRPM0r1xz5yv4+S72rallJvUftc5ddCulnP3Ro+BHD4rU+Gb0dTgXS2IKAw0vo
U5OparWO+uXbZFqJR4V5FjlILVPrM3sI8kMmdWl56S1o48IJOmFlSQjO0CvL7wcg
UxKgNDIXzib3pUB3r+bkyw==
`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`protect key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`protect key_block
hhX+1PRcu8AM31rbT0YGftaKYfcqPVxPmQGeGwpz4LG4g8atkFLzHKN81Y3JGA5m
qdmHkJjn7Rn/PBaAAP0x0siZwIV3Nz/B8rw30HKK8OWpA0yG33GekB4vZlIDOen+
qUwz44lcQbm2GGk+5V7mAKltNSwUqaAZQSXTJ6V7e04=
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 64, bytes = 4480)
`protect data_block
NWVMQzZxbDZ1Y1dvYzg3crTToKm+H0eN7HkK3xdc1lCAwa8vms/JFkWbiyC7Qstp
ZcIYZ5ubnC39jyUxU1FabX5CG49+ZT8KAg7HnTuDVcM1M8Uj6XbqZvWJ/fiUTLmL
I780mHqpJRHYAbve3N8xlQ4rUEQsT1qqePUGcdQ3ONJNxFIhGTiaBmBOe/arNikD
HITcn0ReEKY8VoHd2UYAjLfJhphURp9OcW+XV3T30WWoTfhXKyHBg9LW5wcx0mRb
CXZhnFTNW9Bt2TkJawULk1GyCKofreqv7uwHmFtRhtvJBGDwcbosg4/9oEzMndlt
O8etdrK9jhDR4goUjYPIWvzqyIg8ptaUDxgGClFA15OBgS2yR9sGHbTP+KoYMXkM
FTylPYSY86hcLyjhYamRY0TZw96DMpqm97+cNiLhmEpY1rmiqsma+UpZ0BtUWXHa
4YejGnfindOD3AJ9/EMo/JqrvLuXD+C40FI6UHWAazvZ2peZBTjQykWl4FuZVJPe
w1hIWtJ3LlIBl4Qx78U/QY5scioJmJNnsuj39u+wMIvNZcg8ghd3s3jzgjkBt5M1
stumHeSg0SPXSLAqjsLjCW0MAC8F41FR2od7iIopr0SpQ+D2deX0b4M2MLR4N8WN
QIln7rMNvL4aoOkjDyeDT/0wiSJs3bxmk3WrFwpTMVsHLhTPGBxKd4XRzn3C4onR
GJYZb5+qeExbQ0FVXLi0rmwJkUTJxSGWo1MlApj2u8cEB7C0DImrjq0WgqKpqYKa
BJ15NOdHKiZ+Rf+XjGaD9Az2M/tGjJzINUNvoOaCmKBp0JB3CAD0uaSjIhc8cZoN
QFDovvOM2NkHKgYf3Ws6w7KENU0vqk0YLnDYLU0JoIRNwYCzJqbxFXlwwR5Zxyso
DNtml7NLkQJXK/evHBNSJBP97q3AZ/4V1wNgxMct742Xvl1iEbsq1a6czm3+JN1C
8FcQQEwwkl04kN6bpJsTLh04kjYGN79baSoEX/enHe2ZcPqbMNBvbRUIQcruD6rX
1pKYZ/qKvXlMYP0p/sltvn7i+fs6xvEAAUQ5S1lsSNlP7UczZ+z+74FD7rsgvHak
TqXB8+DMtrOzA7RPsYMvKOTQknaeictzRi93CHek+9zMHvIkkxw2ZvEaY/F3EPuH
PGyFOvoafqgnb2IQdSitSG6E4Q222dRhVPvdT5faKt6BwRamgLGaRwAaR1D5nqvY
L6a+Z4OmAkJkc+HwjRbR7AGfaKeIymnit2qGMSvga+40nf4rdoqsOwtkR9Pq0kkr
jxcPqpx+GQx+rSMCCYRydsXlcBjk72wtu56sFBzyb3yluTXPp2zFPVnC5OvRpGKr
mSS5OEKsyma2h6nkHS1S/pawAm4OAFUtwcAku1WWPkfkLCVoHvH3MUz5ZeY2ZfQw
Am0kdTbjpMWrujsb2dOHyzex4Y//yDLA2DrStdbXJ5fV6UYBWqylOaTi+Gj2rEon
6CuXYPVQqQ6VmaiqgbRT0i5XNug070uq0XLwm9zmZKHaxOQgA/rHwp7T2yFnIX2z
BtDuUE/Guc6uKSmgQdaIZGL7BtnhdoCr9FS5Oi1nZloR2wGlKFq+KDZ0nrdZ9qxM
Tl9EMlJIHM1+P+cfKHeLZHsi9FKTmoA3l3b3UYifGgEUG3fMUI6S/C9pVP8ilaLd
atPKWQ2f0SSVXYUv1EjTX2C3TT8tGOcsdsT+ON9qhWc8VJ+YdmQbajdTWNwD7YNl
yxWpH6RgHRiJhTm5kEjPDjeJyZLAhGo4QT4nlFHQ756NU1usRYhYbl+PZe5SUKKi
O7uuteurb9w5BkeuKnvryldZ67zf1ld8GTcWSZi0GAC06zCE6IPM1pG2kLzS2Vpy
Cil4bivxg1bbfImdOHrJx69p3LFQIiQ3NG9K648/r4Ca6rodPY2OzHTpQ7/ErZjT
cL5SbFdnLZxEzL7e9HMJf9yN6F0+4LrFkWDW7XJmk4muF3dfMkXWACYasy9XQAf3
phYVneUmY5Qy+QnMjdqn4Qftx2a/ggYWWwK9F4+2jqWFdWPA3kA36b7STbcx4x7P
UMqHQmI2Wn+6bpIt6Uu7jw1CU7aIIBesFrr6MDENHdFuQ84etEPMVIVmN5ztpRuf
QTK3/bN5LEZUYdrCbb1lydNr/pYNua4N+cuVakb26YCJAA5/pbr2+quZx40fK8sD
jvd9UP6PFNh1QOYt7jSVhZGs25Vg7fiFlnQlVY5g6/+2CEFOjIjnnUogtnOUPkjI
kdHXxHCZtkdSdiQ3loeVXLVkLS+0yE8ivTzIKJUnuUsSPbb8X7I0AYVil/TqG1K7
UX0sb6DcOG6t1nEVy2sv6zDf7A2jg5DIAd5NxuO+xI0saFmY0/Fu5mrhltfQBab7
FbMjrKDrIjLaYBJpGYYY4VHXPlfc01Ht6ozg4tcVgg6bakwwcBdCRBsqXjtHFZgO
/VFOJ8DLNyFnle4JMnnAfdv0r7WklmyH6hXyxX+KtlXJzN24oGz+ECihI2Gk6hdO
rkiZ9GXZDk+iOcDJs/9Y/jN4fr7TfoOTQ/fJ0zdKL0nYuVOTglyL1wCrycKFtzkG
zBsonno8i0KeYbTG9hIDDRqkCPogCXat2v2n2tmCkIycRnE+8AxCb4j3M6flzGS+
YLE7CmZtofBMWH/snK5dGcxkCNCxMdeVmRzI25sJTOu3WvXhHfW1/jNwNuxsppMa
u8zulIq8X+oV8WbmK/mFH7nYx/4VLHC95GWP3T1riDuFJ4bkE4OfTUpzxNJaMF2c
e/pNj/x5yI1pv1Vi/4DOVTCFdtfoLn+qlC7O0QHwLFzosaoZHw+il79BeQgmM36h
zG16973TWk30Yyelj/f3Rz3kskK/mCVqaoJ3Ot/UrJ8oKY98MAQht49XPegoL5Zx
01a2FmCllj+qVHquEZ7to4kePUTEXwXkQNMRIsHxRKnwcSKkrXZlfRmviGzmhACk
pTzlNr8+UbX4xlGrmexPeVmFSq72cGeEVe/UW29+VTNqzO7CIV3jXaXw9RPDklZy
kjOq6eZbheFuYSzp9y3yVaF9xvaUa8h1FAKi/oDvmrgi0OLFMh2yPX3ZvVa6Q6D4
gcNp2Z9W7Pwwm+S4RGoDAGZPMMj45mv0+N2TyxySwCq3FFDP21xUXnOefgT9jGaO
sGiEW334EPHikrBxYas2zurJa8ZKKdHSSb7oj9QwU5haNRNd72mAS7cHIXjY0vtB
wkjjPeYIhDkGrp8WQ1SXE5ddfRdeDOsxw1eKIeRLAGUyjkQ/EDhFicL6+FnbWeSX
+cOYjUJUlNd6hO+MpuQ85ht3RsZtwVUzv4b+Oiw3OGaum1NR5Lu3f9vSApozV/bp
H+qBuKl4GdDWdc1o89L4h4DMjRXYvkcCG2ibLf+lB5OVoNk2asSarNUCzPUlK2tY
mUJ8eZzsXQZVrbiSnEhXKPgsl3C5RptoRjzeUK9UP91E1YZI/fHkX5uH0TrzKZ/V
aLXNpCTS/CMjPvSoepavoNFLRJr1/nKRQ7orICA2jhqSOh7gQ6XjpQXojj7LxLXV
maVLbsvBscNPXTwE4bnXvFqnCH8LCL7QvRD1nOikOmygLtX+ecXziV4b4cuVmItN
ZhfwllDEj4PV9DNy7rl7dhETKnaiXbmV8NVteSqLbU5YiIHDZ2FJjLJV3/gD3Wvn
kYtd1w0IKaaPu5XSJMejRCU+UAiK7dbPO9F1bFK/R02HpM4Jb1UGjoHwZz5p/Rrq
0rIwlqV4YzKBOt+iJweLk04lNnOf7ByFLMOJWVMvLbLmZWtf3/eMzH/J9awidLRe
fsHqZpwN9iH8vGH+nAlo2kQXUNrJlGtGNr/D3MrY16xEcxYJehy+vZgrFfi1J/rb
YrhvNNXekAlo9WMNdt7NfSopZNBLDI5fpPnvps4vawgmL6O/Qx21YpaEbREjbT2E
akRKkDgZM78NM8pMSxCGextVs3Qh6liRrVMsIHhGeeqLYeUiYev0wclNDoo8bx+l
HQd+n/x6DfnapQZWODB69VTmwJkTAwKuAvj6B5/V1MNwd5WAeqcDoRR1k3QwZMNx
+aQtIkRNHgNEMob7VdKety1vyENZuQzfH6fTDCOA/31js4strlRzl+hmmggzc6wu
xsaETDUCprylRwUgzAUakOIe+Oi0lifUHRKJmdLcagJq27H+CRUJ3HMNRLwUBQYY
pzhGPyhgs6t7eomz4bHpMUcWIl58IypomWe3cFufqa8fOtghwN7ulSIQZi0DQcj3
I3kbRB9eBL5l2oxtiUS8N9LhO9c645iCSj1HUUW1W5WxrfrMkyCsSpLJuKzuw/k3
BS6VLOryHjvYMC1Oc4ybN8iz/G4UisUjJE/BVLBq0TcISPiluegh2aPg8IQFOdVb
KtYgbvMEOD4WchcEGY2IygGAllmr2vQgS6ebbB4BjhqWghvTmzowVOBXAO0pAdeN
at06PtTaF3kiYbsAmABmdV0LIpWvlvXIi3EDoOdn/aqFDEpNi+c0nZkW5CIQOb7q
JY2qFmkFiVa1XDmf96z5tEkPhufX70TFzBs1yU4wEk7Sxkpo93gPbOEG3V5TIHxl
Vkagemv3oIoCueYqgGr11f+OAn2nI/wQrFuS01e6QueugBDLhdqBNMTPEeQkWdFA
hQy5+jnQOCnWXbB4ZyhMWqY4W/tV+G0Mrae+psir62Q/DOsYy3m75CMVPbIYkjN2
2oTpMDt8Q9cgiHKdjacDhnkH316faHEUKRxtunEZTOMxLdDQ5Q/qmw38aT0dsMts
SybyrHGRhCWGgn7YkWHhpFg9XOikknJTqMJKfweb33PZxhb9s7RUER+NwcJj+/x4
YedjbRVgzyRxQJChxUf7Fwr5ajetZj1CV2cT63PzErufXeUbENu/cO1uhkghzyy9
J89kz4litwfO3HGb9hS2CBjot7E+U9dpIDFqdmpFKPJKtJE4GirGM5bljlNVjbxO
i/8yDpbktW/coIZxc+wC+sJAlD/OdLdXx0gVglYzlqeQq+xwZD7yxf5PFasNK/iV
Ofi34YRyF2SjjNdSQnEHOkgBU0azN6N/XNE9qw/s+DkVdUkvxlNWNIPa+6+Ei1vQ
5HfONDimV7ETCSYHg5//ZL6NZjAHCBXtf/OnAAbgcpT4C65jEBHgIHUgDg0T8ayz
f3hOmUfku/odPQkdiybyg+Dn7ROq+Dl858M2dWinj9J5PuWxkQ0jfEcl85piDw4L
htvN66+rjDHIdRrQPYrDoc6zw3Wbs+PVJC4SFoAI1i/8wZn1luDNlR982V1n0DxV
tVbCF0Ez0G/5abPU5UFAYEdNGYVInUXXiH0zQGFtMMqH6OgswCbJut5iFQAMFC97
F5hWQfnOgWg4xQDv5poTVdV5V3QxSpzyZUX7JQgmjDltQQmXer25/443tX6F8fsV
btZyWc9WFeAvrCe7VC1kz1mWn5kY8uceNe1WJ0I7XGD/Twahnw6CbUro007WD0yK
lstrCzkx7SS+HgJtL3Pz3+XdqPQtcqgHz3c647gZkZMf63gj0lX2PwQloOcl23xg
0v3ygv4w/VFzwlfNJ+rQ5yfzxS+rhZZR2kOJny0HzDGwxlTwDDic1NZFWK92kpis
g+h7eN62jEqcLmVyhTChZhhKrowKa/oTtySOI+cgDXUkLblHtMpUP57cOfaKHrS7
lQA4lCa8CVTl+XFf3FQIT227IutUBPHGdvybsRAxDGoHsuHnV8G9Od8xLSSAVp4v
DlRS+4YkRkC4U6/OKc2IpUu2h0CZIHxyPVm3yY2B2zL0D0ROdJo16tMLdocrHQI4
r86CPX0tMozWHMkbMTrSUSV59Gg4uV7tWpaUruBIIj/LXW7wOQ86IJuFX4LQ8ORx
ZjYBBanEL1FjDR83XgK1d+/ais8u5HHdi96rdu/hl95JCTec1lypwhPbawd357FR
n3GDpWi7qfc+AS6bm0MEpPpW74MqvfcTXypLRGi4doIQKKtHAUvplF0NDbgR8T55
Znk74iRUjVWstBEkYkxubQ==
`protect end_protected
